`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect begin_commonblock
`pragma protect control error_handling="delegated"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner="Xilinx", key_method="rsa", key_keyname="xilinx_2015_12", key_block
urVYMXjLs1tcDaDDTEHUqCrcbjaLqxeRRSMiCh1fnAv631K6nOj0Uvn+af4zIUQR0nuxDZLGO5UR
u1llcSNO8qVMjs8B5M5zFRASqmICbZj1FFTOFAmsGkM7UCn062QQ2tBYXI7qUhq0VXurhmscVTdX
ICTIYqVZpZqXd4M86OXw3nSVdZlLSoMiDCGbairdXJs9kgG4oWouCBqqn2XvBrnNTxZ5QPcgj5dW
CaH/SPnYhMZ+TOO6dmjSM+LZZbukCpjezUs1ttgrk+n/A6QjZGyW98AP7ZDrQGRcNBYC9ZR2ycOg
z6QPHADXEblHpX63c5WFMj5CiC5PWuMZKb6D7A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="JEXws9vNL7XMc1vVrG4Us4bsrmjKq32Wkzc+QoSASpk="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22816)
`pragma protect data_block
zDZVAoEYKVe1oaS5WwG70EEDhliAGrjMi8CP74tUvDCWzqdUKbknpRfXmdcDd3getuduzalZGkbr
4p5cuExAZjMMvM2Yd5GyIF81gFw8gF8f9lWyphI0frz4tmtdw1UT/nL4+fwCsAbOOWgiVBLeN+WA
kD1AGktudq4mSM9GKUYHs/bkeLoJbsAgbWSKhsv+P4cdGsXVc5WbNuKXDESyA8SpCANS1725Di6U
HVtjEkb/3h20Jq3ik61+6Okr64XRze03z3MRWtrjffQy1kv0IfV/1xca8gpyUjO1QITsXm73VUqe
OOMEzCizI47weONQu3Ofg/7GCc3ztTvvM0dlyAv9xm+gzPbOoRVFsfMQPB9QczhtXEBj30kaXBnu
B8NcJS1T37IjbGJaDwJwKSjfB8dHoNyGRbWPEgr/Kaea0/w1APmOZzYTZYoS3z32O8l7pziqXZFv
ACgKE45r1VnZK3OIg4AxULpY51WnW3lqIZMzgplEJYvc8JS4pWVQs5lQz/lBk34KEhMXJRZFqd6n
OGLUC04/iJHZJeEEziTSoOejqkvd3WGP+kM2spPHhVuWbPTeb7zH547Wr0WdwuaQT+PWAsZZqsam
wZAIAm120WbNk65ULP1Nok/jPiN/W5ZQu6CeHkY+2ie9OVk1ebKasE7/SLiCkv5rBld3CauwujaZ
UED6VgznFcORHWywZGEyo/WYhZJDxkJXT38pZFjtFfl093qvGvJ3RMSifTDbt0mvOjF1PUv7WycM
maG6r4Fsp86LL59YrtR7TumQU4k9L2J82djhM5wQCLAXArO+6F9ZYyv52x++7FOIP+dY6oq9Mgob
CzwnTOAKm2wLekRVeHk+lWAPKaxGMk+qsdjEKhTLLgC90ywm+x5TU844CDe34SSmaIq57DqhRANo
B8JQgDznElZrv2Me9ZHy21OVip8Jpiodd3hsjIuSuzMWGWMD2z6MDQFlCE03uGFl8JyOqh26eAsI
btuMYxiUxBXCYhnSjSjNsUNwbUk+FhzIqI+v45PY9x5rUohmI5Rdej+yl2tfhiER2XFCmS/CJ2iQ
Ne3IYWHfjeBPaUm9BRXdDqPyhiSYw7BJqDAde67LZfhJcNIAI/CiJmmbBK+ML8E/tzKro7gfDmJb
7YxMJ4KPUU92Jnl+SiPZez9V+FGBGSC5PnmFgotLCl9GyK8/exB/3yswOoCZV68IT3GA5XQQMbhQ
w6fsuAtsjJGukSdhc0wilzSuETcu2dmcGZ/EL28mO4XkWrTkubnAOOEABKLppsQrCbzw7c6valHO
FOOt8Wem0axShvjU9+J+4j9PMwjGaKArd+8AfVRIFlys0PxCEdsJ4yjQwUftsTyBOSZEkAgR3pdG
73KENuY/gWemH9/Jdao3IhhC7RebpnbAiORpETQAqo5kqmi/+/5ixtV7tCbqOL3zSrXyVA6WAmom
bqJ4I5AKSuzTu2CY0wgOLCVpT4GXAQLdusjSxDdZbTImjFkRP5oGVPp8PDWUR20iO2Zz+0A4mLqs
5SS6QZANozqkgJK9qJj6wAOo63M0l7tUF7FR4Cl7uhtqH4VcZaZClxtCgErj/vxIOTyR4+mmnACC
qr4U8SZEloLUgK4GB6VBc/iCAswlfu9yl2uOi7pUe2sJN4Vta3yjVuTG3Gd6Yi0b+tGn8RZEA4HM
8FbvZxzkkfciWp5jdE/AR6avB2tNJ/34B0gMZiEEHeO7j6XSbTiDL2RJo+xno2cwjRLX2Lz4mKj3
BAEUny0hAzUcSMfJPyhEjn3zAbMqAs6QmW0DgdzUTWYsn5M4zh+GKFccuo5sU8f4kEs9Kug/yC2w
jy2qBFIddpr/ylbPXWSAusW/I5OZqaEnAdTJk8h5wtXwbpJvZ5u0HZBOcG5N4QY9uu6CurBZ74Ip
dNIQN6VpbQ2F8+Sqhj2+HNWVwRCX6Q3fOLiSrVnnVP8Y/dC6CtY8JjpQRzPKz1hmQHraiCuRiLEe
1BUxr+1ioxVl0D5b+UmwbVwHJVHDjfHJI75HzASgyk5n8Se484Na/1v5PDwytZJGy/HaNhN5nYd5
mjGGirbUu9nAH8ayQRYSHLTquYHffa7b1l2aLS2ZVD1BPjfpTnvaj0dMMWYc2jex9gFOc3lc0jqO
NWeOjNkZB6JPK8XbvQJ8Jl7sD4D47FziFlL+5SrVUmJHW1nftefHT97Vr7K/Fd64CSGNq/sPKAjo
yQWMjiE0MhwbuT+24Q2lmhzHSVuWTeDQez2/jY+5J6i+KWGJlSNNqb4h+oo0cp6YGIGYZqAqMexa
jVFu82YGyxhd6ft0ccu+pz1m+i03YTnsYZIaAt22cZaA1SoLRA8RCZvxLTq9rA1vdDNwFWG5pBf3
Qvjuu4wO55nbVCIrf3W6WWExQurDbs0N6Bff4icoaRUUhS+BDmacW3TnAM+g951TcnYtN4SNLO1d
oa3DcnKu45/HCMTckT7+WS7MV6w4x5b4nuee1WL6aUOfrT5En47+MKZ1+hD/tByN+EEct0L1TGJn
X7QxupqzkYNcGbnFYAxA4q+HHHZgp+Om3+J2KBdvXIT7X3AHRqDvFuB6+6mY0GPBoA6qIJhi6Dyd
7OZBT5VmIFE6KzlAxoIcwrrb49tZJAsVVvihQOXgJfhU5w/7cAr6/xUMLSa2W83VmAA0+CY1hmY4
Jy6SpTxHyCJuDpZwJxhoXRkhwU9Q3oVSPL15ZPJMNRTrxa9wEir2tL8JE/rIkJfZbpBS/RPUuzMW
HOnQ4UvbHdCcEdw6i1lApmgikUfj1VW/ktIsoohe2szRXrLHPFASikNZwa/jhITvbjQWS5zkTw2q
9ZC53Eo3p0/X1S8eobKwE6I41vRgxCc5mXJnON4+0/f8qQmEixx4aL7G/hBFRQNIha+TdkCWU7BC
L6PtTTjCvzlXgbIbk6ZcwJxN9Cg9aKIxTePT0EYznxLtuSRh3YHU/PiRLb+tlH/qJlak0h0FlKc/
KxSSGZDqC8bz0ESq2fPGkR8DNYm4+ALkA5eCmH/4MElTErkUGn5a97rZsnvgvDeC048x9US1Ces/
gMwgQRstZeY1VZRIzuaGxZPwxyovxWFFwo6jB2QArxzk5jomfVIM4W6nCPZedzOAXfJSxXovnZ56
ojQ7zFOUHwnjzkOmEPDB+WSOE9zhEV/yh5c17RljQ0ejBUxqiHN83w26olAvvPR6suctgZ922vPq
GPKLTs1SwUhBGDkOqL3lcslMqdgTwOJagb5Z9jujiQN5pmXnXZcxiFOVPhGYLVLmW1sND+wvOAD4
M6qoRnZ4Y8xKA/OT0dBJx4Lvwgj6omsfe/q7bSM5NamVljA483ua8KuTbwQFPNmNyn12ywCIgTdF
pAjZhAZZiLkR8CA9Rd8s+6B7ZKICBK470l/n3iSpuwTEkIWNsZKl9g6DeNpXbo+hJYF2ZDrv7Z8+
eBdHNcyftphHuiFMOHRKNc+GbzHOAOFKuO5FFz9vdbSgv9IPL7B4gamfB7SKgfh9uYG0E30rRH5Z
VfX6yip2OnRcnch6TB1vZA6DLf+OwLrJCSXx0IHuGkVEEHN3FVPVAbwPp/gzeCgX2WkA7/Jx4dXV
9KWUpnaKvk1aHEDa3gCikq3zgw2TA8A2xwYvRVWQDCkt4kfVnGPS6kmuLojsr4C2vj8QV+7VXZWF
MQnzyJ7MrzIoKY9Xt+7YIzPGwLUCWLflQwZFmY6KKP7s+5ZOwFUMAXRDczc+IGikuCaHWhtl91t7
fxZdsDYcnxOhWiUdvCPKsLLhYyckSbhld8qLcCfNyZiy69MfM1xBkGGhFUnqANTi1FSsK2tNQD9h
WHIJd69RMnKpi9ihwPs3ZhDo32BQAvBp4ibfjpyux0ZjvzTyuyzLZfKY6UlQk9rhDWMbQf0cnDYe
pBG6QuscufMcjA0+5EIzMBs2wEi1QsnOPKAR7Im5Rdb8XlBdV2K6zWGbGrtMFKVBzgyEkrzsDhg5
7XR6DbIR2c8r/xGYKo6WGTi6TxeIPZeGxWheVyu/N7QytCg7keTVybXRRTtEFuRN9CuLStcthMRR
MiV0tBE1PZUJ4va/+E1KUjZ+0qcekvYwROpiWborLCSFp1HcXeA8gLtbrg0xDrMILwB6JX0EU/Ih
6hzu+JUZoGZ3e/iFHToDaqjt5KLzkGkvTDtJcbafH0rgG+MA9f5I0WG8c5SL8LqQxmAv6HB6eA6G
0JZrMsQXbffRQh4tZpSz9IZ33E5Fe3bI7Lp/bp3XsqW++lg2WcldxO/hO4+lzwpSbKyZjw6E0JDv
l1cNYkyBoZjs13+S7otKu5hs+gZwK78SXF1nNZEb1mverVkZ3o+p8Zdp0OEpYwW/gHN1ZKG/31QN
1HriVrhTKTk3I0oR/KKvi3i2alvlvvrTsEwEpjljIDAj63H/x4O/LiCP98ixKSdMg8JTQ1jj/JaE
T6RrlO9qWO//TrcgRsQ9zKNG43Ge4PWvsjDMzuhmyZcTPzpzOhRPgVQHwuUXEM/Tjdt/4tJvWlUv
z5ZpvjglcRqqSnec00N6QMNBpgbGuH97fAh7dvoGT7mRF9rL4EnTelejRu2YI60roCrs/eKOcHJt
8l5wS9zh5F49AFpFcwLueadlaWZCgYmD7E5QtBc4BIVJ7qHpe1sBZ10zMPxCidK3Ktlf388nVsmM
4AYdUwjrhtugtwEYh+fBKO5bZAa4FC0af5Cb9BHMjpPBDXt7LtO0aHxMLZWCgBQ7JADn4tiU0mSH
Yoy7Lb2RmZ8A9EcGuVqEuDUIsFaKyGOjUSTRNyBB2stFMfseJ21n0YCxpR9aFx0y/+XJxaRQe3t1
mB9gaNxVriOb+SxFSiuCxSvrK3jsjJUhmMLkoMLnri9K4+yOurFK7D8z0QktXpwUYDuH8E8CP/kb
1Wui16GdZfdvMupfYR/boz+ogdOChvdZXocxR4zLir18E2XgEOcxkc7/5FEgB1HJ8jKitsggAojX
gd3QfazfVsvnVCDchKhFt3+5fl9TgGs+d1tjzm8pQelAz+vEbHV2M8FG67ZO1p7AJJ7JUr3BKCiI
dfcQAxSoonIxOvfJyJO1HGtbJ9NvWk34AkjBhw2fbA1Jnh8SWtJEW0xwGOAaCJOUz0X6a+S7ZGrq
jm/gbzvxkGQ7xlskXbSUb9VxIc3qJLLsZY6WHCA8r3kmTRdNXIiLiwlH9YJIfKs5zGqZN8sOdMI4
qY5h6jKGlNdvsZ0goxd+LE6y0az/lEYyNY4K3NSyHjYUaXEkXs+vSIH3QCihEVxfN3aTKmb3J7rx
VznCfX/fjspV5BPeV4+RFwT1idV2JFGjakrG6j/LVGG4FPrNUkc9xLnSgfE4ZSjxDoV95Ow+RwCh
FzwiiOJFjuYp1TasOqkBTU57as7U7Ec9vM9EPnoNguoA/dylX4nkoXfghgGlYTe8F8iCABUh5Vly
ISU953IxhAyFWUY0VRBB6O3r+zqEhdzmpQN5avA0f+IFDejB/ajtMN70egquQhUtNPrhyBytw/U+
+frM+ZlEeYT/h9uBkNbw8yGhJBdokGFyUP4pFqut3OsuSP19UmnotkK++HH5jDb7dJraQyeLdYpW
2QTl1QlqSXyx6PicTfcZfn5gLVRuFOKT6VsI6JAhOsLOD6MBiFpjr6Y8qZ5KAUu6jlbCe5K9z7tS
dtsxSff4FVgB5QoXipw2FvBi1rd2nObpP1rTY65qpSehZ/CK/uVg1LYy70z6eRPZH5q4kT+9FX/R
NQ12Pbfr3+193q5UzhQTTdSz8SBtG3lKu9cfxz5bs3+V0jgXOd+jguwIm+tZurxh9AttPzF+NXxC
voH0sq0jzdjYOVFCpQNjQ0zAV/NkbGgoY9NEuHTdQjYHYogj3IgHPjzcdnihBR+R2Cim/P1fp9JH
ABlGwG0t4liTg5VqMwFEtvyWA8aqzbr0jNEXK3TLqK+dEpmrwE/+kNY25c5aQ35lbsC9PGAnV20V
eIix4/43bPq8OsvVD3iG3AWK+YKAbvu9y5IWkqVVWgqsesUQ3hPCEU9JxpIyyL3W5IqTIlimkAXX
LQBTReQ65xnamabrOh3m1ixIxaNNf+9ByNhmfFAy2zMj+QIoB1y8dfKjPn38O3VAJ4lJjvgZsKkh
0f1XYwDM64g/LcgjJefutJnHfHcVHb2dWtKMvwax37zlACszu30gst8CBFNIOb1xR7vMAu2NSpto
7o4aRXUmNaLp0TtC2koQ9j66Eu6++0JzPjDDi/TVOecYkyvgdK9WQDQtWw+bi0rn+jgWLD23SOh7
6Eu/+6e1b8dckppRG8QOvRdBG684G899/unrCeXg3pFF36OI/WTbdO+Xy4m4dMAXCHjhxD+2B+08
dk1kvoz0K1b/xOcJnERbR9ghrsJccJpxUknS9ryAdEm6KbXTGzQ0XWZuqrsGGuvPMFeZDAJs6y+P
2SKUZ8Mw1Ad5f81Vk9JDKTe13vuJP7K9jXu28c7q2Uds6cBe62Lf5ikmtDfMdyoo2rfJNmnK7JDX
6M2rNT3BsGiVNw+WD1QbuVlKOfLBFYnjgTI+IIW5JOc0MkbH31nyrwTll6PGJsNblEIzIxqz0/4S
5WH4Ts1c71R3kP2IygJWmBkzR0bARqowDienXmxoJQ8OJa742+uIbMEnlkXC6ihqHDGoUdHGN1Fn
CwGin0/fmmKYKkrwsyhQ54+hMUqi1LrBH4h9m0aCiy/cAx+pzO/2A8jkK8BMmRbVQmQ+kjNiT9yh
BDXrpLtFIeFKrr+islVDnrQLhvAUCcWMnW5nc2j5LQFyZvPAbv0OfUJOIhMgeqVl/6dwGai09y8s
kte9krhi+8dYFUt3YjnMPtWcDqPxw7YULY/rcphYb+yAtsNF5e3YMy1MVCqE2C+VRSPRTHeU4rq4
3+oYRZ5r/LE1D3TfMAG0YB4STijnEZgQg4zS2oyP41D4WvUtQwlfDcAEsSrWtlJK6pOSig6XhuEk
GweniG/Ob77HJK6yFi3lAiONpqxuk5h1UrNkbwtCLKEVP9DyqWjlK9diZoHr585dhwpBcsWp4wla
lVizhp1jd/80Ct7lvc6rEfe8GOULo48OUPl+xEtMww32JmH/q1oJ4ho2bMHFQN40fKXWLfiidywC
oCcHnSd9gdowQmyuTjx4a9j2SZ8sFukrokWkWgHxOjbpGYE8jozxJRwjf6vbbDWirIFVRxcq7P66
b1WjjmLN9GVNfql7xg6DVgUdxxHtKhr0d1Xn2bz921yTs1H4s+vhxkkudkcltqH2r+HcNYXlTuLa
m++Zq+MPsTw032UhlOGzVIaXGM+eeYX1ogDeKYMm6DxCity8JQ4qHuYcY/vCY25thccimpWw2Is5
Za40zBJeeme2DonlqqTcAf8GF/OsBRz7bQmbOwvuHsyqie/SbLm2SpMu1P3hMpo+EkbJ6lZfAPjB
6T92z8frkrGsB+E4fVoTjGQu3qdxXYx4B/MYjQG08UD/gB1OOnBBjF4FvGGfpLMasMJDTU58o44Y
RJZz5JFWwK8DJ4WGlkDnDZmsJUB5+txsHSGkv3C+Ioqow6DQSXKP+Afof5tg7+oF8wGDkmfvqT3E
2/wFCHJPD2frZe4tPDrrpj9On69XtJElE8dpy4lUkB5NjHNchT6zWAHojgRZ/P5w1577QAB8bvJu
1EhFvTu+BkrRf6336mCboJfjX/CbypEAE1wNGAQ6LAeX72LMpDmRoLVUmfeSNlMZFxtenmFrEKPn
7QWUv1unEBj11aHcyZm//O5S4xZJQic7JePOEkcSqod9ly+//VknSoMIGEUU+4t8n8qoYVL6Utbb
qCzV3qoS7lxyiFKw12C6wru1GlEXnsYYzHSl2zcdgCbbX/kMv1TYU1hnsEehzqr9hL1jeWZwQeha
3oA6c19iYy4xuveyEYs/g30dPzRtPG+OpH5cqHbnsfFz4DZnSnm+XRl9Id0gcdzkDOxml9Dk4YG5
1InwHgNSSXPutGBHN9Iu++IMXigS8lATBjF4747/PkoiZ45fUurfNBKmvAJ1lSswRZTqwme1mJXA
EmsKbgBGWOJLxcwwEqG5j7ggqd8mQm2k9y2phHa+o1ZppNYoMwYLi3m034Lk3/4mV3SIv1F+/+5u
/AL5EEMmt4mS2jUNLl2lE9JmT0ZxldFakJ7SFSpsdl0rD8VfJ7lZYl838CUfHRk2+rCBE1EZ308j
Cqt3XH/XbwJ/+bBdkAfK/dZNc5JysZcV78myFQosfwVlE6KGo6408IG3EOodQxMcWB3ri3xfpf0M
GDhTWlL/5XyGWsZnsT16l3k1vgSpACZkozmYIjEi/TWwUpDVT7hRgcbQU0waHFn0XdTE34YORK7/
UrIGwy/DDoukxZMXTw15UjymE6aVEnrKM7sY9xE+A1TLYmwkpFNKtZ6REGVZLNbG/ArNZufqLWPN
1M+Wcz9SlRFLA4iBmFrXwzqitCel5TM38mzNgAulVDpiHuHAmdQElkqs7GxpaeKcEl4WwA2MPeaQ
2D82PrkgSO/vprSwVzHpJPcK1An8h7rUwI27kfPLT16ju11VDkWrujH7GRwOLDYtVzwClqDrROB5
Np7D81oVweOV9RLT580zyI7jBpqTMDx+YibMm2RPgXbv95SLWk8meWufSYdCygM3FS443T+MCAvL
pt9G+rcazLujnLvpHvHjT9WfEQxhA5Lkth+OVl0dDPRaNh1HJ/nuwuW6rCGFSGmxta1cpWi7/g/E
mLvIgb1umGh71X/ZsJt7shSfnd7hSnf4sTRIHKI8UQO9I64w9rrbCyik/Y+vqPCOr0mcJ1lSYYhs
rH3miGl1ExlXsnXFLviz82y0OqTgSJVwmgEw99XgPK8pahyzf2Hrol3jbMQiscnqgOJudNVRDKze
2CEOApeZezzKGSGzW6Wzx9qv8daNWa6SvemQZc8cH0DN8zkePAgthOFmEu3rwqtjfJGCG0R2vina
XqQhC4gTxXAlmEH7HwUFjV+qbXm7WDxuyumzXVtNbDsUHsB/HAZ27bX+mjZqyfZotUEQff+EHh5G
WVqBQq2UMiKnPtKJGBCk5dM1W8AZZl6gL3S9FSyw9c/IWBScfJI46wy+ap6TMICYPKX5DvFPR9Ww
Y5is1iXPvISQ1fszyyZSJH4Sz0XG5YXaLQZLLzSgc44JRB566kQaqaGFAd/abPEYkmwEu30h8gJx
9QLAzhCyjQOsBg27X/FnN0ChAsJBoG9luttOgp4kwD6Le7cRRdAk7m0OBAJPT4Xj6kY8v0IDkU3z
MDB1U7dYP8sL/2nS5KBTXKvDEXdTNdR8kimIWfXrPZfDXu3TBspKF/1Bm0J/AOexRdefiivxF/nM
ZndMljyCz/0hvc45mWVAbyrO39rcDwHXed82lh83leieYitOlnUOo69eLYiYw7wF+ZjKDE4xIV9i
f63rfirj9yHfA0znkRIUxTVCYKxs3PxfGihrQqqnkMcPcddk20oDvjbnVnXP15YKoAFp651N5cf3
vRoG6/MrgsLR9kV9vbEzwTwxcqsIeLLmNviq04MKDkUABSNUg9I+fxP8MzUV6kYOq5K9A8UgNM2x
fh5SaPoOvr7w2SgcJx/RNSnIjsTAlSHkhdYW7VkfelCUxYitvLUxsp9+QIyf6K5AoKSBlSMLaKxB
IDscyVgda2mzo/bn4CivOdcD7hD3SR2S9jbwLTlqs29yjn4TjujoEGRQsBZDtEBuzKgELB0tJHya
GP0syuvmV5Ebpyc4K/A2xTWzqeQUiv+Am1HvpHA8usQ7dNTsRaRBJlZwS8VUK6+q93emLaaSbxxl
pfmkeIW4XSuVQMgiei1mdmmz30p7iWEIaboIAUkJZyn3/5ssRamPtqScIEo1P6V2JLZE7FNaeeoc
d6RUEBqossdgQ8cy2oWTGBBgITq5UctCU0cbPT/ST8qW1ke6NhVvAEtT7MvWMJHiXsbnl4+t1jUJ
AOlOjOi7hStKraGiqEc9FQLW7eifddMkUwEa2QtXAgFMrVyo35xnN5mhGT2ZTBZrwFHEwZCrYELj
JHod9HMHM8OQR460vd99bpjchxPdlDOqa4DFgCMPTjjPzGBwxKHRI6nTamP1CjekJqaUb/hRSpbV
n+5PMkY71ahFKmZVsn2xGjpn2IIfkxCbBtjBHqYqtNQCfWZTIr/P26/WHYoHk1ITiyAXMPhmOIO/
4qEz7cgucj//d+79+Vj6W9/v6+iaw3FQr970hYssH2jQgZaVug2yvGfP7MCsZ59ANR/uVPc8haT6
rjWZHk55fbPtNvx6vNXYQwHCe/Q05G7m7/D0RFtWFOqcUf+8dL6Uxo9IbPh1yKzOhNRCCvZZQNMF
E6eKD72FVICY7TfbDWax60KnVWFBbc17p3XtJVaZMqoUcNahWHgMcRcE7/G03Z4nJGL3r2NwW19U
qQrK2HxzbKP90iBNuFxS060RvuUokmaSVez2JpWgwsZ08yQdX+fNBoZxGLFB/lz3cpbu9tYSuOVT
RR+o14mCosNWCJLKDoaHTKU1Xy7IbbrxOgEp7l0I2m+TkdAYcXm2/varSlueWSI3092DdCRZY9Ay
os86bishJoUjW88k29/c64giPELce8BH+x/rvh3HNwnTnSFJxbLJWSOdkv4a8FScVPYIPi6XzOhw
NhEfOmlIgEEASBc3Xk1J1EjsOLs4SGOXXrZxhFnz85mkgunA+B1hvwjwqSxzdZr6KuHKLIlv6XVp
lH7AICvzK1uknwpmKfX6wbENPjw3UGieZD/APP1IUee+PWx8JiwfHTy5juxSui63Y2dGsN6FgO3A
TTkudv0vG0457dCChZJ8Pv3Hsrs+c+Hvpe6nWD9F3iAwgr8gHjbsBwGJh0BdANFZwnVmFSnOREL6
ZqQtPDkllc5cyiBsUYqnqaDXUopsvMSZOSwMmi6lWm0AwFTSUMfBVguHWwSKFObCeiGfm5kyuNvL
jCNCPYOcpi9fcEqs5HYTYniLY9HcC88//o3jpSX96+H1D8aRSsN4RiPLs5QF5Qb/a+pRbRZIV1aO
CVE05hlj/xbgmFLkYgLkdHWHFZ6FyE+WfT/JiyvpHTbjOKogdYzdVffZLhXI1hVbuAezmoSGYx4F
6XZ2L6n+8dVZR4fzVxJBl3//dnONBmXweKIcCrdFeGqLfUPHqZS4hFToKZcorqHfaWSvRe/UEd+V
FPTHV6+fcaERFWPNqrx2m79tzWS+XNm53zjEgUfykMTQ4W5zWUbpcugzgo8l1jsCU+DfS02PP9uD
ppCj9hbQq4kZ/nWwbkOgUuGUd6/DQufSaio0Wh+F0F3FL3Nk34yn1n4msNvhbkP0E72rAFHCihMI
3Afx6vxq09CnezYAtNcK1tMZEINEKJ8NFQ80OhDLCa13/6JVnvqGxItNMiqH2dvFp4dEjvNASkbI
0Fu4Mm+K08wTUYNeawRaK6OG81Enc7XokJVAP+Ozf9xSt/uZoVTj/nSKgd/xMIGoftouRXYsn8FW
FtyxTaOKZvC6lq9tqzs+xsRMT+niX74lNCiHfgHp65NoNKh35axc6j51CBG7fYcYkocOypiIaKLH
oVaa95Cr31BTt6Ly8ABelK0pWPF+b1xE4oMwhuS4+s5+VScPHaBcMEkfUHfgDaUEiLuB2ytUv1jw
9adNz9py1bF1ja/G5pBN/grZyJTJkK9c5ZelTQFttMfpbBksRhY1xdYRBXRvLRjDoeVexMMdauJd
t/n5vdpatwlUerF0ACgEx8+vc4nr5gi9rnl9OiNruQi04T1vggEe7n7nPI2/VlH4InOaGKnxsZsJ
uELjeK+bLSk+pbF2pNcZXhZ3/FjBgBm4Ey5ZK1ZANDwcvOcrxzV9JSReyGmQ8yKQ9/JnjUDHZByc
Vf+4JtzHHYK6ukAthsO8toX3sQEzK62sDsjNcJPgO+buDmhJVLZc+KaUI9ilgBeSoEJGbH1b1rJr
bRcusIN4an62Y2NhC3eHNH86HsJtYcHsYMHZDQ2Iv9TRv2LZartrll2Xsd8BN4xaB8ZlOr26Gu7X
SWEb+3YBTjJpqX8qCWYhtH5U0nBteHlKOqNYZuz4Y5+t8ZiPep7l9K9lavWSaWDkeHZ0O6A6kmjv
eM1HChTLIiewh0vLavJiPb3rhkP191ejMO1H714GIISo+rWs4+EsedLRwle5RrmU8qbcJBWZOMx2
/+1XreWzoJVmXiH3K804fqKwX7nA9uT/ESKCFegFaeE4N34g83By5V8nsZBlU2faWZ3aKBFFXkc5
7Be4+vnEN56eJYkp/NmKbC1c9zkErwEZtv7PE1scEtbNqlhu0mf0+oijDfkDa5VcKb69jmYpSSru
XMW3W62Q3tLtKNxJCFeCJ1PoPf0FN8bpRJNWx/0umJPm898rTMApWfb16jv3IQXszh0vifXOQ24t
8P7xKIisyja+dG4t3v6vH+hi/3XH5bqNL3ntEg/ZW5gcQpBZ1wDDvVvwduFIW0XDZ+8/AcvTYvVH
nJ6JiyL6gFUrIPOePiV/YqAdDOChbZgK3nM2PuUcTtAP4zuL/0GVsDdMRi87+x1URJPyGMaRzohr
8LjQWsEYlILJUwZvDzOxhK0VAfJRWtQ7l/FFW2QJty5HxGaCOgNCFbVxBWqe2S+XMIuT8kTvIMN5
8CiYBv1CpG3h6FSmUEw6Y1wfMfCE/dKfIc0jYu9voK0bTMadWgOpozvYfXh3tXCG6zoyrR5LlVIo
adqAKZnxTeeN9OXkeFKR2CBe0n8/ewHJ4PKWx+TtbteX3TfC+sNvIi2olcVmNEXg2gjEnlKtwcf3
6XalzrfKSr8G3XaL947hrxfklqdGlcJIKHiD1zMYRGOBZlQgOTjohAHeEW2RU3xiYToqsQE+sw+6
T/1OlOddVTPj9mi0BvCoA/e0okodfKd4SbMFVjHvZLacC9f2o52AENZTSDEgLD+JtcPoLpYshSRp
rhEfngvswzUhfAZ4P9bZqwx0FELReB9K+AkjBENRdXwnde8Bm04LLQ6gAceZpUXU57b1H5beMR5Y
D9TF4XyKuAOuhiAZAGf+it/VJlvphQss/66bc027BpAhPV2pErWjbAvwrV7GUjobWgrpRWc1JfAP
4ObhBKfjIkl0zvdzaPbwy9N9gLWk/jWy71XcejiwH0E0tAuxHh9fN3a76i1F0ENO63Gw/v9Z+YFx
X8sL+vuL/lDnOjRgZbQky+rESNA+RH4k5l3sOIZo0M6x/IuKhvtvgqxld4XeTPEMLqmA38mG4APS
UdtecWKDAhVvC5dpa3YELogh43QGhQ0P2dF/BM1E4xAfiQTVdwRGTW1ci8KJ8U/3DklsjOuhr8d+
TKSLep7dZ/Z2u4x++C5YcSiTFevC6T0g0UEN/Ik1KZP0WVXpXA0GsCmZAYfc1f2ouHzagDoNuZAF
LQUNUnUekR28mxDdck+uozfd4BQ2oR5vmMqSL76RYKqLO1X3HWFeifkyQppIA6pXqaq0x7Hc1D/c
aZm3aKyqqCTWby74bDlIO0uyrkqTHKtGZ9lFSILa7I5bZQ0eil52b3hkGDC0v9iK86ckfkk0lJig
LrXvDdqPPjIXjsmNdNLijmlk7YXLEIiIghnizIIYbfEccpDhB3U18kjsZcSp4697jIUiFvRYdVd0
382D3Rdg33tM7GWHEsdn+TyGLe+ejOplAWVodMRJ6vVoK7/UzfJ1aNuJcTfjcusv5VISjrnD1SBd
c1RnWhRC0mSE2f2qv19dEPGaRpgcvjPHtIVNKWLyCx2UrbYEFGcs7RvgtO3H24DumJQfK/mfM/OX
8Hhzj2xxfH+qBbVRfkI4b6l2urmQBeqJ+STT5QHLLnyBUPRKZPPNXjdJLqk+Zs86/HXTEXiEKsEG
HFPF27/2FhhCEBsVnt5LvLmkCLe2C7/rJ9K3ITi7E0zhSRiPXCxBqffqGY5yBx2IOy3bbOUQmpWK
1fQ0PQlw/cN2AkRadKXDkHcupJAy+JK9Cjk76sUelLobcJv0t1TMp+1AePiT92lBl+/F8pVTO+41
/U+UzllsSDqU67aDstApdnzbp2LW51cMqMfImOc/BHTln43UAC6IQaMKiZnS7eNDgcAfqCM5likd
6m9FSpH+WFVYjW8xVM7ImQt0PaEKV1bxQhfDs4X/rQzFlbe9baSbXDqLu/w0dPdVEhnywgtZFMdz
zNBzT66SC4x9bSr29ppVTceBVZoKkujMZiVWTTz8txLcII0uz3M/7MBQIyrQzStb5s9Z64gUonNk
IApFVdexUqSYRyfcU+Jg+DaF/jgh6wnGbufJPMM5ku+smyBxxIP6ugbMwPBfaTMC6qk0VliphiPO
8ERJQY7cZJ7DCzSGuMs15CwUHTTXjg650nzwq+981P0aA1SFvUYL7M97s6lVo1hy7Nzgn35BQTzD
JOZVPHdVyWwbpZsaRt/khYS1noW/OarlrveR5hf3+iRUEQKZ6f/PTH0NoEMqZvUfQgUVX7i4wQFw
z75N91N+TipVFOHXwH5uTw5xvNg7+7mkkaPIei6a/ByfXXv/5uYa2E2NR5Kwwf1UXmfrTisRp8cp
eDZtweAL+TBwJg7DYN2QSs5+E20EIcr94uSf7MgRmzpS3EZ1wSBBG55OZutT+0LYJf0xEAAEHOh0
ZQfFdZQ8dHD6qCQTwMPLaN4RFxjTD3gVBhL2UxsGM67IUtP3z564EYlgKlC4WioBEuhdKIiljmMP
r+/67Uu0ZNQuITPj6VGnBqbjl8g35SBcIsrl7/u4BNh1dV3wsuB0WivHbpx0uGFoRXq7vrU+pxlI
iXs50lTDXz+OY6hMQ0C468PA5uIDsoyQwa1TnnAi2JXO9UqX/91bgi9Ozulh1NxexF3LlH6KEtUQ
A/QFgJYuO+70/U1NVrZ5oI/c26bqZE7WliXrZ//AYN6TIp0O4Lw6BDSwmOHbkxm1Le3LjGy/Qmuy
XX7C4C4eBcyqGF9nmf2HUpXcso7VC+eB/IYeCEOGGXROHOjXQrZUbl6zvjNrk7N+EBFa+F9YTrwL
AUoTsm6qKHe1J8hnxDiWJBIieSIFSzN/rlbFC52P/0YF5HuKr74sZsPkiP4rYB8BAKt8ytsUJMtv
0F6gAT8+QijFzj8I/Gyom6lLreMJQM42d3NE5Wjv2p1qf87PbpzYlt0V6Fzp0jvhrwPvoeFgJ9x3
Ei9eJP0nk100rAJ7Y5T5F0gGfGc8Qn3ovXHwnYp9wlJxYlIjrcAc3YXaOmNL8VqTnLx+hq53m27N
KAB5+RS4dDcZwVY4ZRn+nBamgcuVtt8i0lLQrB1gvdNNW4+tibtFTFLpSijiPWILbv9LiAA5rzO5
wb6dJLbX4X7kCBfycTmDXfKXyi7a8BIOBfJWsFO9N//KYJWFGqpa4OI/+2H7HRk7HILbxr+scyc6
Ib9AH+0TUZ/nyv6sKzx4Zo7QGu0EeIDsyTEmBFMDqadEIs0OgNVDKSFDM4EPIXHmpkxgZGT4n2GA
tzD+AV8caGYrR09+nErSfebJZBUdLWvZcPFtVqHWcvhrv8s/1/h1fRthgjrU1PV46Vprqlg48Qe4
pLKPwhbS7fpbTfOx7j9JhcYLpsAFGACvERZDyXWKNJMJ3eqsuE96Nx7IYBCckpyncLi1ykxrDAKP
5BYU89k15UgzaRNEeaeSy8j2q6b15qSX6bgxKKiAaaWP4rGohY8BWQ3R1H9JiQZc7jzpXbQtElJs
CU0+b9nU1w6CoSbXUrl4EfMt+fxj2kvw6qA2os5/UqTGPeWoPU5hV1JR283O/WzmUwlfZR0kPp5r
ZnN5F/G+7pvEfLlfW20ZWbVRp8vbLveJxZ06l6ZwFFZY1Vxft7/GMzuvF9xPN1n7SaWT6kW5XdDC
tapkbTSefj2NgAGgk07Tq9A1+9TuZbu/Upz4nPKmM8oObR3wKr6ixQQVYedmuMSzzPJRJE5Yn96q
xWf2Y2DtxYO/atvfhYeV5AxXG0MlToOOvM4umJaQqGQR2ZbuaYy5kW5n8qiflBJAZ96NJtYFwtvN
IQBUptqM3HWKQCAwJZYy/QirOtMDCU4e1BI4cVDvqYkXiajqLPLJ6YxchbrvIJ7sZAyKk4m1BnKu
tLC9VwvSkLy/jn0cv9DV0VKLaNVXk7CeL4HXMAWRoO+7MGNMd9xwZta2cMGq2IpS+t+uHlPzCHBr
wU9gdSiMQdd/MZtOXqEJWBVV/d1hZCIPFAddy1YnHjkSGTSDgTsD6/8ll8ZAXLTb8Bh7SZQ+2T+H
9kI8PdGV2QnVVgiYaflkX6M8Nhgmy1b0qDywtDw+MzIc6e6s9j6x2ThHlkG9OMd3ujJAJeXpGEpw
cNpAN7vT8zth6PfTnCIRqQSgmPTV/BV8Kl17iNx1iQ0q5EQFT3wqq4n1Pda9MPkHMPDHvjovJXjn
jiabtc39lk66+tni/JduTQDNzAwcjVbBarXKEEIQYFnkaJtP9sPZJ6lZMTOgDT1d4U2vISgEf9DI
3h9UhPGbQTOMsn9T1IHSpg/etsMVk2awlsZGKSfrWbGoJFGWqZJy1fNzmhkJUJg2sB/jxDgO5M7C
dyMTRJVeAiDqrb0+RWzP+aEC6UNyK9n5PunUlyw9XGgG7LT5mSWPAemYVA9Qcq1ZnQjV7VRywF1j
0FkjGF5k6mLal0spb7hqMchNjm1CrwFg8LV7ZhUkJ1DAvfNxZfXpGcyzV76QF45HuIWSGgLGTGAj
aUQc+8bzzdCNHsRJfEGUpS58DsR+FAI+rxtEAd6rPI3g4jbFSyyaqNP3lUqVSISwTmljnDfwGtQj
LgTQ3D48nwe3FTowcfhMuRVRdLuZtKQC3DKT5T7sIIvbTlRbCqnDDgov94iKLM3OFRPcmmUhw0yz
9v6gdhp/v5bz32vhmxaPBLTBIvWCLdLkjkknTm8oVWUpXjnPIp9nrPMO8JxZMnaENsmWLbKEKyAo
0+dfnw1KLSDRBtOZhSoZwcPF5xpwh0KNsAsn8uB0kmblnHFY+5V1m4KLCR3ZUYqv66Gv9G2RYLWG
4+cLo34g2KxvRfXCyzUilSxyaca0dqdXgjf8cY+Hs/Ci1RoZj5EiUSLQPzToXbL3u9F80RLncOhw
eXO2tSAS6L0eAOU0EAIQu233Pw/N+v0x9FdCD4NihaLyE/7CWE3/OBdXtcjoyBGRDkul5BPgfYHL
wqVPYIihsLhNqrn9HyAX8dPyYGfEYrpgLsqvpRD4Xpdu/mq9pprFyHTMWBwB3Yw4AWyf0aT9qXyH
zh6XrMVNQKTkuw7svfgqAR17MRzmuVbrTa7rSIy7dll0U+iutNgwO7LWMBR+pO5V3L3jSZQOVLw5
bqkino4tbMCJ7Cf/RsVGEPGAPh6FtBJNDVN+Ida9LHvsurbCaoPT+paTwE82Q9CyWhzrKRHq14iu
hRzSKi+FHeMiUdoTEwMSOt6yu5AjuPivNbbtAdLbpctNZWVFbu9Rcn7SxhyliYNlxiD8BU5vBDKP
7Mf6u8whEuhiRHTihCNuEK9VDbODhmYkd6jFU3R2dFwXaR4QMV/O0snDh+CNnRO6FozzsAUnPtOb
j/32sveT1EX5USfJgTYivXLs+NksgpsgVCsxUjJAPA5kc9coCb+gegXhtFXgs/KUq2E39UkLpuh5
IRuy/XC5GFjJBIej6kr9CxU9QmL0ICY7vCPXza2pIKKSIqhJeQcpIwAZN0U4mtIW7Zu+5bD/BZpE
kcnoG4A86GxCdH3DvioJSTV4mlypxyzQcK9OK6bd9mSHEDTK0PBTNxh/iWVcvotevEXobQi72h8a
dVNRIyj+L18OiIkqSh+N0IacP+4nPnLMeoQRhtol/1spolNf+eHOG1EOJm6EBfpkEdx2tm8gokgf
8mooZJE8y7XEQvxhlqVcf0tJUoKwD5nRHJ3LTg3rqPGDO8EmiiryI1VaZiXsbEYyfzqNFnbxYQFQ
lWTXg7orPbthcagCg+BYg3zBW/I5gVsZ1wVotGXTt5InIQtBlHvkKkUPJaFIdDe9uxQHjHdnxu6g
RplxjyhVe2PM+xwJorjKdsVaukxJtxWg5iDjVsffKoHhWLZbD8rlwSz3rGT60RhLI8bBis4v09Gh
6ROeP5Wdc5Mbgz5JEw01PHCVRJ5ddrxw9Oyw2va9FP4AakhbNyxcdyCLSUmWo8rEppjxWbhYOQoc
0jvgGp/O9XzKsjgKzTr1cI9IspHfiFI+TpbmzLwCTYwYHjwAoJrqLzDO0dqrsM/+F0g3tvWe2RXh
uye8jR1lBSgQE3/QFb+nZK0oQwVdTokV8BWTlz/8rk6NFI5e+9wmvDhN4KPnhw62XNvZhJqIlcpH
0fg9fCVZs/kNbuqknRK3mCyZ33eswtKa3A+/jqR4ZMY+8X9zXfGa8rLV6Wj00Q3/MB3W/czb9hNh
A+YRNFQ2/XAr1r50zDyijtQMUqRC3B+RBITj+kAtnintt1RIZMO/WpeZlAM9RwcChAOMkdZMoi/L
pAOfAz1VaVkfZ4AflOXFF9lj7Zexgdf98OoVeKA7nJbxxNjqG8o0MFDNvTy9wZShbwHF1c3l76ot
cl+r9n5Kx9OIFaJ4T3aOzqv7WAlx0B8zaXGNEf0orW7eVvcqKUnmuvz+H+uPrM7P3XhUvJmglRpR
WVapvRZsAWTIvKPJEFl4bDLdzfJBE/JPbQc2f5YxXlMKX8Eix9fjbYZe7lg3/fnqX9ioM35/akq1
6IYB/hjGGRURMzaIiNtOPrfBR6FHaJB/k8OChuLHm8UKSc30KYXqI8zCMnwDKhp6R+UUP8AgtBUf
kvel4FastbD8rlXc5CEVsrOG7RqZZXxn5tllC+7ZSg2oJk72uWN/LiI2b5Fj5wHbjRLRC4w+s7G5
gtBmr3JPg9NAZ8OtScjdFB3IO6vP5C2jjmoFgUGI/5oml6GviIZuWiHS3J/uNKJbBwuR5OqYEG9H
PLtp/4UKaShyPfw26ZsC3U/n/DOT7a7mN+VhpY65Pv5T3VRWlmTVX8K/YwdddN9RWIPTyBoclToq
/yB/pyCVVxpZSTxsajVDjXiVSmPa9lbh7q+KbW5fdO0EqojqGxzSq+WXOG32OqD3V3gHSbHy2Qsw
/a6suVVQavVmOncGO9RpHZ9mAOj+zbW2YOiFMYlCpHl47iVPuJZ+3UcrdvvmlnzPD/zLuIyMlTeJ
jbk8Ik7ZZpg/tM5Hwbehd7KF6rKrpNt30ez/vJJnzz6vX5g3XG6eDLpAcRE5KcCSJOxgSGmLm55R
SjkW8fAQ49TH6hfX0I2c0qijQRrmfVwncRU6yX+jZwIfXAcRGecr4qRQ+LsHs7NVRax3KIm9Gmj8
i8L9ogCQgNRHGn5A5TotTtAM7nEq008kZmqk7YfjJKWd0BS+7AZnRtSDA4hIcBAXkIXnjyTTQx31
Dk9/aXcSUD9YtubXJ2hHjE6bQb0e6A8twWAULxwDrkk75VAoqG+fhfOILPB6wcyEPGHA07RKf5tE
S25Od02u/BfOPiY/wtUWIdJt7aRlxCo87qPjMhtC9Mjqmg7ZppNIx+oFnVGysUP4Iw68T7x2Se+r
JnlyI5xTIPJmo+GnkiPQNmjD4nYDjpNsVqvv7kfIu3phUY099UA0K4lQczD4we3yOHSCPfr1Xz7y
2ly0RYGPqhH/3dJIsPQYVG+6FR1f7yw+wU0NH0YT/A86Hc9IWe6sEuRTomap8YaADHm34+1DrZr9
tsZ8NX1ThcCybveerSiVvL7wW+NkwRkA27gglPmyYJc+RmsWSsveCYdn/5hs6d4MuX9r2o4BJkao
uKYfuTtV+yuF+0MrysTcyjXVh9uxzlWhn4s3+lb+5XwnLeOr68PktFYNrkHrzcycyhWkiB7pFr+J
l9kjk6DrK4ZQqJoSUuYqCCI8u3vtsljsg5WvuDcltdmg8RSQNtoP/aXgS8do2Ly5fce70fxfKyt6
SrCkxwTo0cMyhuI/Ntq2g+cP/RBRC8pxME5i6zsqMDYrBfCDc35kbUpObA8jSsQDb8BWFL9GJJgX
O1wSfWU5JAVAtZfWi+iMWoQwWIeFxLtR+nCEGyQoZLoTtXJ4yW79TZGxspTS4rKrlR87F3nDz00d
P6vo5WyVp/y+Gg/GrViNVhEdGmONMrePQnyuaDdK04bGMQM0MtErLX4GmbdOYTVzQVHbUUsSmU5r
hkW8sN9zsbzjrQT0e9pYewT1P8Q7szPt+ONFwRusRdS2y+UQV0W/v7+5FIHgLRi1Y4pgiCpXrh26
DMpKurgOycVj2aLenOqAOgGqrLfIlggAeKmuF4FLY25EXasW4pXcJ3TiqZIgoGJgJqMWoq2j8HPE
EViOEQd3K1xtinr+XATV32SupNJ/Q9l7TkZsjff+5KNhD9Rxzftbo8+LRgC+cVzL5cRZawKmVmC4
fa9TMwgV2ezH0oaa6wwXYc7d4zmzI+ApqtJpEofwmpwttW6Kv1mgfIN+Kn0I38t4qTNJRJmtuO6w
uwVWT0/iLnvevHbzAD/a7lXssyhrpTG1759B3bmflRjtWSx0gyFHjv7UFYpbVoHrHzXVLErleRtF
Jh/ffqijQw6Alw8YNv4+IAzvXrWG4fPfPN/f/2Ew9Iy5s288GVmE1UAGQYJCTEPFAI7zHKLxghF6
+LJb9YxpC3PAzNThrXAUYk1RRdgdCc17heh1sFxbc2/NqR98oyKFLjqMMptbNrriF0abIX7iUDEP
VXo1znuR+KtxtsjDmW5KpJyImkqdBvxta7dhxqVi6d6xTtSIL7qE3LJPJeugQpdEo9CHO2y639CH
bytWkYyo+N4nBTCrm4yT4hIdRjsZ4qWqgoTuOQe4+JYGYTTThwzMvVzzY3EdsMyHoZ00sOVLvCAm
n26DeieiRjMOcRdyyOQXua+v2/WlNyx42XAtW2c6YpugtgXxogQ/U61F0bVn9Ofjy2aFy1KqeX3y
EMPoVpxNylePMIM9eO7hAvYWRR3Q6kkksX7gdG6KP0DlE393kHPtH/k0UtY2L4TI8cI4FKFnCmPZ
u2p9355xz0R9h9I884hCangISFOnjxqt6lwY5ojxljDwH5IfwBaBvjjAF4s2dRTWVfxyTkEwjPfu
j4O457pYUBWg6TJIzCQovOmYuny/uldtoYgVM61q99orhC6VplGSkib+oOY2AjsetIUMTbKkC0aj
P/S96V4Y01pkE94Ws1MbQGSERIhgFjKwX/jel9n7ayTjaEUh8CFcuGB/C5rToSVsohkiUY1cw5ar
yQK35B5WZfVatfHuRF3EUHn91qe8ASeSH9Tfl7cZzWSNDIWRdf9PmtuC6FvavSRteMYITw9U4dCq
Bwcc4zR8N6klvRVtGsn1ilQLXzsfYM0PbI4xHzGDoEBzqWqxl2TK3ARN+Cqhcj9rkppcUn++GaCl
hR9NmYeCa4Y/6eSSnUFaMucAydQnrB1tbZnWgJesjomIXom5kX8azHZ8qYB+jF2DolCFqER0nYZa
rfQJRtb54IGa6PbpVnRtio2wWpTMxy5LiXjnnCJlPc1o8mxHsHsnPFo+y2Y3i94Cb5ZYz5+Utqyj
ygJ1GhrPAqkz1eFsLyOX6LtvoiwE8oVJ1m49tETnaIUJYYZTlAfYUY7INsx71bt9Gc3bnZGqrNtA
fowHebIZ5DX9VYv43ZdIZOxDpHiPY18/tFjCEd/OQj9xkwjxrgAFGtC8YMMroCtzsN7ubR8ZOv33
i07OFdfflbk2DNFoWgik6G+I7yxpruPRaHHcVREyRdVL3uL2mbyDoXTSYh0p0x2aGCutGkgCB9J6
swdh8eAQd6wwzWCWj2zFUxLArafiFFfQmOPvA3xnGn4rAMlR4q8w/Wn3KUGf1hKc6kubbugDgaFM
irZwDHmzgLLk5pyaZzr69T0cbzThvDAo4iwqxeujPrlGhqjP6cwqg3ERmjYsMhlRwtisJkGFA4/3
ZkAh1gik3WA9l2Oq1O+AYWbdOAfAdnKbHbYu5Ebl+EeWXiUCrLJoad67A93DZtsPdPpW20lxBgmB
LqwrKxCX20LEuK/S6kjqkauoqyZmYP4DCKOK6SMUf4g6WGciJZOuHwjCjPVkDf2MFe9bcmD9lJBt
zz5PSGK5CG3pIcK7KAKcWiJ7cwOWuMI2NaSvqGtaQU7RIuR2lDOB7dhngOQiY/GDtjZU5LM9fufM
xiPWy/4qiS/nQc8WKx66RqqMeIHM1F4E4iesmSiSh49vvgVY0rHUDgb9w9pFN0XOzWc1PvhocFs7
3N/uq9iY+B/rmuzEW4Ec0xs/eVxJNLsv7Zl/Y6NAWTPdF9N4i32dHyaT6+C4tniiXMN9nPvN3TqR
YNiLVrw5KwZq3o2s9O5QR36XbVRtypXtVMUMxJAnBYQDWqDZw81lFm2gkpSYB1bKWQmYvxyYOi4Q
oZO/u3crCpKBs9kbwYpS5w67iBLLCdUbElmifzYPgmFuJ7sTOopPN+r7qIl/APy/tVaceEp7YjnB
ImViz2FSPp6ZA+DL9uDd8LxoahKsuTv4Yl8rAVP5QdUJrt0SPONu7qC/GQp0TO2kiqHiiLM7R12f
hiRaRHyHbnwJMzN2mtB0PIeYfpplxkz/ajJnAYwQy9+ECmWLhIoxau8PvM3w7IMhXo6KgNNwX8NH
/JOSo4d0PynexUUhDfgGHq1YcPPFZwJbvrXfTPXaTXT8F7F1/S+IQA0Xg3uKAk+kQ3kaX91cKipI
dszdYORFrUE8i6gKx1IXrjuZV3eLexbi50oJOVvmtMOb126hMB9NDHbsUvXcsQgJw/dAFIzwnapf
Nh+xbUvMgan4eYt7Dxx3WZ51adgD0A/XuYQTF7Gv65mkYxGPPeQAd8xC+cuMUFzFZ8GsQrY8KR4T
XUGUMLXmXC4IPRzDzUmiExp50tDemCixF70nW4AwL0ytlJBW67b3MRswVrAmyoDgJ+Q+RobjjD9w
VSXF6oUA5RWSb9Z/XEp4hrj0EWwCh528rCmRFQQ8TaSix86MkSVbdHY72dftfuNfPWVrhi6DCSE2
L0l9FjbK+gY05JAKMsAz/YgXkOfIOPHZnAbmwcuszkn8/5J9D4BZBA2jpG6fUgEp8JTpW5oWjkVz
fgj0zlKX5MDjAhU27vIBG3EyP1wOhGC+Y2Wvb2gG2nRPQQT0j7EFXsi8s0lFQYjMZNxdo7ZDq9O8
WiqxBKiBpqYjWOIweal7uA5fPFsfrZJhHIaNiJjW2VME38+GklxrY5EZnw9kpHzRaoJzigZQzy8T
kRhRcPXGd2MqKSbgzEBDAo0LFWnOEn5DdxkhLC983H5h7xrq8AQ0V8o8dpCG2pkK1J6IoHJiOcQB
Z0qkARLm3AUdxmvNrk+JPUEXqPfg2kpiPz6AIZZwNQ5rJXxldCVNcNMA2o70cH2quKDl1G5QlFLN
WeB/X93XqodTcJaEMLCClda7+HRu9Vcn4fgwWELiIcKDWxz8p7HqdTTsPFH3qnbUVcvbjaeQWipF
h4BLR2N/HVM9mVC6oJVCaDh926QpuVmSlyR5hXdWVasU208jQN1za6BtcFsA4MF3FCnntzKy/xlH
2J3R3VH1CDCgVAjqtG2LTbmE82+VF7EeSbOxV5G3WaIO//5xtyXl/WqVcrHPP2/O3/bxmwMUmAKz
cD3fIr+g3otgGmA1uDBwHpS9rUDv5LdAKWdlzEQAfFHDmmwrCI+cVpVVTzPFAgC3ujpUDvVl9Y8z
xfYykxX8QuDEnV4tbMXTO9HY81TgKAGEogeS6nT01zBnfybJ/RagD/PNZMCNzEaE/a5FwRwVtAyj
IZsUWBt2JKDsbAr8rJK4nTf8vztlBjHyAxrKenwiuLpijo+9K+vZ4R2LhkiqZHYegCVZPVtsSXT3
5tF7HdXII2a95jXl/vQA9IDEd4w8Kef+cUXAdw7pcl8u1GntDi4CsslxuiDC0kMkmmYF8MiJYjQd
ITnnqUubGyLCwkhtBAsmiU2cFOBgghed7IX3RYImV93JrmkJOkP/GQqgoKBAR/7xtO4/7wlP8aqH
CHE71K7V1dreom9deVy5016r2Fxw9co6rcmQOL7rFCTjlsYv2GUT8ok2XOXfVVDJiY+G81ep68wm
I9Vtf+yLY2zF0U8JgiBzc6ylLC6MnGIbou+2XGmDWVz+Av7T/3aQSKSz73+qgodybs352OC00arW
6Ipg4AZoo2ZJYhuhJ7+o+/rv0B8hJPUmSM8MclnD2GTzKc7l27qOdTrfuIFV0tbC7h1MhJc85VoY
inp2k3BMU15oK9U2djwCj/ZiqhZ9k8zxn6/g+iHDDpt6R/I7EurRnxfVKVGus+U8sHaJY/O1PqsX
YuKit6Ja/d08SJjMYFuXKCuZ4YfzhLV58e0/7LRBTAI4Wsnj7MFvKTCTv2a57Ng/9+9EjbrLKOfC
uL4F4KmkDBCLbb8Cb5GK7Hb1dCkO3ifcnJS0qrpwZpQbMah5+IVX0ejVB+5YNhnsc4Lg2DCmkGgL
usOnI1bzF3MMU+fu+COGGtcBL63dFF/Mpd6/aPyg4ksRkMl8kT/HV9GjLgDemV2ayyNsh89xtxS1
mUf7GPUUs+Y6GHzdAL0XZSwRMWR/stmJl9KDvl95kLNlXLGID1M7gogTGcy94bhQ8EFtZm7Fu5yZ
/+45rnKrB3eqmo4DsJqk2YPWkHdWqSj1Kxv90u5dJdknIfJkSbzVsq0N9N0wBIEy9FOZ/QjNZ7GF
ib2cjnUhUWv9VwWY4PWwv0yDiPdR/wzQ6n5IkoBLd8dREV2TX3rkN83O3a64e8NoZHWWctoI8ttG
XvngLbZr8OPwMT9TuBqnU7ZMytEQGrbMkIEElW0537tPxn6W157fAGV9Z0Nov9stF2itYYOUXTTb
xAZ02Nv/AZUl3qRBd9xW6whwWFKwpyaZnuKywkoVBjqDswFoqbTO+PE+T8AGQfZ9CCQjnsEy4i49
RiZMB53H1GVfdXVr0q0ZneXruLbSXUSRTuykXzTxdeX9F/8VA+YkcY1o6TDRYrJddZ/pDhz4BaNC
hTElJlFBdkv/3lCKz7zMUt4uqd2/jdR77MWdJN90oSq0ec7N6mRm4n/G3NIQe9Ru7xbTLNIJvlK1
ln/Oyu0n4SjV08iC+80Cv6Z7b05jhx8u+sbEhxPD1FMOaOIr4Gq65fLuiH7Y5yr95pVRtLiBxyJt
I/Eccht3vw4u84D3e339NEtRojYUqLuXfbH2ynfcmfGJWLZS2Cqg6yYZgt6AJLkAoG14PAY+FKlQ
Bd8RpbTH3BgejzR8A5tMvksyVyID0WlfjmEYyxj5voPIYmFl7QBnjj/+dJVAXTRlJic+1V65l+Ao
3mbfSdnixx51yxgVkxDfQQNQo7bIee7TV45XOLxASLq9/Qd1i2ylTBHawqmo5lEo7TXbHutdxqpn
KWm+XnNfbqwHgDc5jTsGsVC/WQavtH7kfODH8UBAsSDhq4HvASecKsFjm1Rj1QPFsAirLi/p8kck
L5zaJrL2cxwYFTzl9Pqun+Ys48Fmmm7N3YJKPC1fN0b/X0Ux4IYVES+EOlJbnX8DcGGoTVidYBib
XZQi5+oo+J7sGJhlk8vxjW6QkI8+bv9UydLGbCrMiV0xQT+nKa6eGjlHB812HNZcD3Y3dJSCcg1w
7KPfs0ufaaoyjii/TpY1AKGI/yBx7rlTf1X3qIMYAUSeDzIWxpw+l4Lr6cTX1Vfyj0lynEy+IMvs
sRiRoAnutn4GJCsIOS42sd7O/T4Cpexb7OfXfv0Mn47n+BrJzHoTis6HJ2OJV6qF7DZ5wMTGkXPA
Mbc5cANR5P8IZRAdBlHpLx/OsQ4G3d93qHJkvxyNbdwHqrdNzXBQPuObbbgLgZ6ySa6rXTAaPq9L
Bfdedpr6lWxfvxXUkQSx3N3hZI01ED2xq3okpii5vG0pyVnmG0ciXtArnoS4GSfiJuXRILGbeXKJ
YXTcG6bj5PXDkITH6o61hPg7LWQbgq7D3H/D6N2+VPrq6vTzqfPcNOhsZklx5CCbPX8ALD1mstG8
lAfUbEvatktLJu8qUHwIbSarSNLcoP3FI0tkauLx7L/Bg79Mgf5nGb95O/zKq18WTZWj8xRUG2Dh
YGWsbJddTLgxi6XwckEOK3e4GDVpw+S6zrQxyzqPtPtWiDwQy5MsJt8X99UxMkHlsfvNxbzjGHbY
7srAOT9IGzBGRxmlUil/GRLWyH5dHua3ifcfNpuUlaNN9RKEuv0I6xL3TaGFR0aLFK2DZtVF42kX
0IHRAWYCHmXPGxQKd3YTGz1MOrb0Vv76SlB+nlerUHvBM58NJnbgeQckvo2iqcMWLGY5D5frddOx
WZp034qdMa1zAgoDzVp4EMNxzWjKubxASXLLVMkncUplZx/RLcq3+PwlzcREPADp01b1ZXXCYz1e
t7YKrC+vsDeG0dGl8n6iYpCl2Qc8rHJJx6hYt+jbB1jME8SB8EsyRQNXQ1jLpUNBg9ez7JyYBT2X
Zn70u+vOEJhkGcPEGQkTdwL8tY/M5tYLI2dbzOlKqBOKOodhdpRCXnXJIC+BT+8AzTRzbwwhAhPT
x4ACBgTvXxUWQFBd+psK8Vs2HjqhHiOyS8I36LRwuGSTufuiQVyKMuad3cQCc81QdgpUSo3ERs9x
5oRK+6rTmdZ/k1fkqcBr3MxpJEpYUM8RqZtb68A/P8Mts8HE9Xm85aspqPHG4NDnn7sLrBcPb+xb
aJLFZ5TbEX4fWmjfdH3QAgz8CIVBg+D2MQD+GH7F5vcAlHOULJeuMxzbOreETmybFEftaIJlERMr
cEggpyQh0PvWTeZXLs3y8jqhimF6fCeZte0gmWf8CxJmyHfSVlEZVp7bcQq1GnA2wF+j2IRFR3ai
Wkeyww1ED9XneGnfYzCteyrxYsk19xAnStQASR+ewluVj8i94kfxDISd9m2kjYoLhCdZ6/R+D/9q
zj1caEkiJR9kXiXSUQttIoxDtEJqJt5oSFQB2/0cEO6qlc2IKvtbH3CbWhpkjTDupQa9eOYlX/SB
Fw/ZD4pvsbv2ODbbfoewvqsLON1t2EjBV5LjeqTSWj5ozqU0HG33xm2saE6+VO6aozCf0j2Mqhse
5i3TLD1RtCJFweO/AKa77eyDP5gQWwifgD1jLD9QKDbpraw9A59OjuJXjOuV2XrQOqyInW23Ma1J
L8kZG7V7XagDr5EWpXJ3Obww289nXpZbpnMGASLTfpV51zPrxfVXrK1D7WQznlILVvAWg7NhOr1N
j9XVK9CfrVwmdxpWnmrqyzxb2xZMThj54L6YNpr15zUHlLp0yXTWDLcfBQFIm5cCbVb+0pHUMoTx
aDvDqhD2k7Y9oowhyOYpaKa6usATwyp0eVBIhrfnnwOPTn9DdPOrxry8FZu21t9PVZxTsY4oyDmf
wiTXz0ziqtsIVegpUf1Ki1sduG9bSf2TxDJjU2gzDaU6Ifx3/3kLyQRETAauYONS9Zc/nGRJNvwf
Z5kWOh7crSN0QHcDQ1hYXu3lmjrZeXJLemEioJA7I5EInvqQB1S2zo4rMk/8m6oXAqOJYZbZ8DyM
t5Ivrv6IeGqneH9XU2sC7lmEDM5AQ1mmbWNzZuGuEoWe/t19/uyXdTN+7xsm0Lmxpx7zUwU590aW
i07/DmYXAadfDSzciZYwtmKeULU3jblLYQKZVei19iaIaa4qPIn7supOHnTONrJecRItXFJIFspw
UCmYiYIBEEElJMpCFJvooeb/EUhGIJvmbQL5y0zjy0VQRq46TeXNRxwc46BaRIjmdKJ23XUlzgEB
BBL59yLr2+6dINUDVott2ck+meJvUK5mCqPWELyD2E9+XLOnkck6QJpIAGJOkp7cmzyvmS7ZyPGP
Z50F7jT2tjFhIqLsnFmZXspLJg0OfP7uerRYd3PFe0/ez2b4R5w4Rm6RZh9F+gLRiBUOwVD7fV6u
l499btb3MEymbP77MK1oyikos2LeaGsNOxw1lA8ZoTKb/q2JMhp0RwgyQLXIg8TUfPreHuaJwa2B
0unWRtvl2jfH2vfCupqO7hQNctjb4UquQnt5ie3Hlo+PJ6aNN0ajyHmi+2FbKxSENK9noCh/t6zE
sfs/fJaZRu4FZDz1DeIlYRmSmXGx7DlprYp2QWEt96ri4lOcuOD0NTwFwOCw8R8iyQmWol3E7Mau
HWkola2nzxji9/N/Ic/btE28VtJIyw3iIXVWVjfFTu0j6PD77KQ8I1+uci9kKRVHm3qLsWsioe+9
4geEATiAtXolNfwLlQi9HMuoEak6eig0HvpzQccRl/F6HOq/eosYP5sD1qGvhsVFeMIq3DUdkaph
RKH7JUx4MCsF1hqNuqr+0R53BWhgZdPxnEX4xhGfBs60+8LGPyMdOP2FpReOydn12Uw62W2hKBLn
nNqxvcOXZSd3guCi53fZ5evAkh7+BN6acNuDmTN1LC1aKkBsrnQY8PU/Io7PLpinSKE8vbzVu7j5
M3nR6IhNz4afQWOhs8C22buW2B09Olqk/pPC2gWmh8ajbtcCaqsbdwFJAc4hrLrC4oXf+URITArP
yutXIouSrI2851wsWADPAFPY1uK18nx83aRh3QSDyIXY/TuBwXTXC7uFAB2CBej/M9u5XQ6kCKEi
xldK8B2ghI8dWkegWl0KU3oSYgelXA8P8+sQptb5MCctWeF/VoN2/kHHFOkSYWp98LE2mkmeykGm
ox6M/9vqa1iWnmdlBqECxQ9IfghhPll9XWMYcQIUQUUGhs1ULoQN6Vb1o8wV816AYSi1A6XnJvU6
J1JlCLOBTJso06TMJ09MOUuY4K8JBFvdrEcBJVZvc/bgO59X9l7gAG6BdtpNnWwfM+avAYzL/Cle
LX+VmF1Mv/FWmYfP0+YU9IQT+eSOL+lDUGGuMGRbiODpkxlvvRCqK9PWJ4w0LhYzqy81pNAItb/e
3Yt2n+7wFzGUoUQZ5uLs4/YAnfCVfxC8aFdz5jK3L/7X4Z4gnHbA9VbYsrUKvPfoPlOZkD7t1Mvw
OY4zEMbc6oQbhmoyNX98YFyWZAwsrs/NmwOlg4JeljU2a9kJD8uTef66J642O75V27ZHLjnAimDH
pqDLGU74EmbplJ1Cxh/0qyC/oaHepNgSYgX4bNUfV4SbSW0n7u0w/UqaacUwNZ1V8uCPDBpn+dWq
sg0PCVXT4LIUQ6Z/sDU8yNiga42iKjALQZh6+D629VGDvc1Tl32swBqu+G7byubBiXJia5JF3kd4
gWsQk8UJ+B+kCrfVo0rwOaX1ETXkMXXBj+Ffh5VYrOi1iSWgKWOG+vO5Vsi0kaX/HUNcZW1UZgBd
8ObL+qdNLt1MgH8+AuED6TH4/zbF/f6AHHtuzIMtbwbKh4j/1UC6HyVa33dJKFCyIL2/s0//Q28U
GrSW0RxeJPEhiC7Q40v8jUztWyd1VT8tU9v35YXroARgaZvBGQM0mT50B7+RV6p3V/DgRMvy+iys
PjxnUoL6NW7apSfNTOhSV3nJg5e87lJuC6Mt7ZidTJrKW2J3VEvB3gnaV34quDJVLlfImpZ3oW88
6xlsrUULuuZ9vfrAOcTqkAVZAWvhgJq2/aTAzvu+ljjoIfJQsvNmXigwkK9PH8+T2+dM2JrLjRIq
OokDR6ipsqc7j+A4vDdOUmtmtQTzWkeCR5lgYWxf3uXATHqjirheYf5lJiu5b35zqZ0XIPJ0tcEr
9Gls9n5oM+dzU0GBTngM1fGJTHF9s5WmGrHQ33eb9PhdLllrHpSKJb48KjIw3CM8oUYs4oj6Ix4i
uVfUdNIH0DTCHp8X5vTPl0Tzw4uJj7vX5HkLzXZ/eJ0gh5EsO2Xe12Gy5YTOZjO9U8MMEPHgl+Yd
I8xypxv/JXNHZC6w0UxsQOVZZDIiVdQonfBwRK0Cr/e50KXQMCqSgE3zUtx3ChlL2+jq/AZaNYt5
KGuYV+Y2u0KXDSozie2NGjGp5QT7/7ps/Vy8dO79dF9RzMK1yztDKu/R2O8i4pRO7omyCMG7gTBF
M9zPp3D/i6m+0M3LWgqZbbmpX0NuD2OUhkzNQobPhwfrUnh3f5VBzzViwSHGQWRlW1cAQD7iWFro
NX0IYn3/eNr0drFXIz5eHkkuR6MQzc9BMLRKLL47pg5jKb40verp7uW/7SwFXF0ryGbeCGYEU6Bt
TarxjVc7GHrdKeA3x9O9NNVuDIn4k89JhCjIAnP1xX6BconsRLQavMN6z/qGlOspelaN39iZgaBw
P+R4bvgBZJuad7K621tENWI88PlTyH42Z40h9YP/NeGEuAXwNB4iO1twbO8MT3vMJWpJY10DyA8V
08QlZUcyktuuuUfopyTKdPZOhFHKLWpHjPJpHXQ0F/NIugF/+P77MiuxuteJqskdZmT1uZ5dGJ/d
uD8QbXSkIO7R18Ohg1OyEAWZyGitHNwnA44k3wV0b8oTtvv0Uo9l4i888zKWDrj1AgkSPSb/SjD4
QoqqkcEYS0zOL+qbJcLDxUhxEAQxCPPuxNIFhyxu0CBwSFFF+bTFjhBqHWkPQ9aMZ1OZ9MCAUpcr
sPuo5eXBWlkhXBBgi3BnvEQV9OaF7+lFytC9fcr+eoWK6pkrzrilx8Y57ykcJYAz6vt1kFtMakzC
SVEtLNBinnbLKLuC9od7UBjy2ItRhZbjRuUDPYEWLW2N3fysTCzxRKG7XTz8ymkpfhW6f++lZdNb
eYPk/0xTuuNSnFkntsR09A==
`pragma protect end_protected
